module adder (
    input wire inputA,inputB,
    output wire result
);
assign result = inputA^inputB;    
endmodule