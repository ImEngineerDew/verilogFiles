module firstFile: ();
    initial begin
        $display("Hello world of everyone!");
        $finish; //Stop the message
    end    
endmodule