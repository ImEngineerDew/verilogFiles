//-----------------------------------------------
//This is my first Verilog program
//Design name: firstFile
//File name: firstFile.v
//Function: prints a message
//Coder: imengineerdew
//-----------------------------------------------

module firstFile;

initial
$display("This is my first program in Verilog");
end module