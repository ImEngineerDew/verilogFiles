module firstFile;
    initial begin
        $display("Hello world of everyone");
    end    
endmodule